`define DELAY 30
module or_32b_tb();

reg [31:0] i0, i1;

wire [31:0] result;

or_32b or_g(i0, i1, result);

initial begin

i0 = 32'b00000000000000000000000000000000;    
i1 = 32'b11111111111111111111111111111111; 
#`DELAY; 

i0 = 32'b00000111110000011110000011100111;    
i1 = 32'b10000000000100000100001100001000; 
#`DELAY; 

i0 = 32'b00000000000000010001010001000001; 	     
i1 = 32'b00010000000010111110111111101111;
#`DELAY; 

i0 = 32'b01010100000000000001000000000000; 
i1 = 32'b11100000000000000001111111111111; 
#`DELAY;
end

initial begin
$monitor("time = %1d\ni0 = %32b\ni1 = %32b\nresult = %32b\n", $time, i0, i1, result);
end

endmodule
