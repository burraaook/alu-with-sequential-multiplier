module and_32b(i0, i1, out);
	input [31:0] i0, i1;
	output [31:0] out;
	
	and and1(out[0], i0[0], i1[0]);
	and and2(out[1], i0[1], i1[1]);
	and and3(out[2], i0[2], i1[2]);
	and and4(out[3], i0[3], i1[3]);
	and and5(out[4], i0[4], i1[4]);
	and and6(out[5], i0[5], i1[5]);
	and and7(out[6], i0[6], i1[6]);
	and and8(out[7], i0[7], i1[7]);
	and and9(out[8], i0[8], i1[8]);
	and and10(out[9], i0[9], i1[9]);
	and and11(out[10], i0[10], i1[10]);
	and and12(out[11], i0[11], i1[11]);
	and and13(out[12], i0[12], i1[12]);
	and and14(out[13], i0[13], i1[13]);
	and and15(out[14], i0[14], i1[14]);
	and and16(out[15], i0[15], i1[15]);
	and and17(out[16], i0[16], i1[16]);
	and and18(out[17], i0[17], i1[17]);
	and and19(out[18], i0[18], i1[18]);
	and and20(out[19], i0[19], i1[19]);
	and and21(out[20], i0[20], i1[20]);
	and and22(out[21], i0[21], i1[21]);
	and and23(out[22], i0[22], i1[22]);
	and and24(out[23], i0[23], i1[23]);
	and and25(out[24], i0[24], i1[24]);
	and and26(out[25], i0[25], i1[25]);
	and and27(out[26], i0[26], i1[26]);
	and and28(out[27], i0[27], i1[27]);
	and and29(out[28], i0[28], i1[28]);
	and and30(out[29], i0[29], i1[29]);
	and and31(out[30], i0[30], i1[30]);
	and and32(out[31], i0[31], i1[31]);	

endmodule
