module not_32b(i, out);	
	input [31:0] i;
	output [31:0] out;
	
	not g1(out[0], i[0]);
	not g2(out[1], i[1]);
	not g3(out[2], i[2]);
	not g4(out[3], i[3]);
	not g5(out[4], i[4]);
	not g6(out[5], i[5]);
	not g7(out[6], i[6]);
	not g8(out[7], i[7]);
	not g9(out[8], i[8]);
	not g10(out[9], i[9]);
	not g11(out[10], i[10]);
	not g12(out[11], i[11]);
	not g13(out[12], i[12]);
	not g14(out[13], i[13]);
	not g15(out[14], i[14]);
	not g16(out[15], i[15]);
	not g17(out[16], i[16]);
	not g18(out[17], i[17]);
	not g19(out[18], i[18]);
	not g20(out[19], i[19]);
	not g21(out[20], i[20]);
	not g22(out[21], i[21]);
	not g23(out[22], i[22]);
	not g24(out[23], i[23]);
	not g25(out[24], i[24]);
	not g26(out[25], i[25]);
	not g27(out[26], i[26]);
	not g28(out[27], i[27]);
	not g29(out[28], i[28]);
	not g30(out[29], i[29]);
	not g31(out[30], i[30]);
	not g32(out[31], i[31]);

endmodule